lpm_counter6_inst : lpm_counter6 PORT MAP (
		aload	 => aload_sig,
		clock	 => clock_sig,
		cnt_en	 => cnt_en_sig,
		data	 => data_sig,
		q	 => q_sig
	);

lpm_decode7_inst : lpm_decode7 PORT MAP (
		data	 => data_sig,
		eq0	 => eq0_sig,
		eq1	 => eq1_sig,
		eq2	 => eq2_sig,
		eq3	 => eq3_sig
	);

lpm_mux7_inst : lpm_mux7 PORT MAP (
		data0x	 => data0x_sig,
		data1x	 => data1x_sig,
		data2x	 => data2x_sig,
		data3x	 => data3x_sig,
		data4x	 => data4x_sig,
		data5x	 => data5x_sig,
		data6x	 => data6x_sig,
		data7x	 => data7x_sig,
		sel	 => sel_sig,
		result	 => result_sig
	);

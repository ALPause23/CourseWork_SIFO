lpm_compare2_inst : lpm_compare2 PORT MAP (
		dataa	 => dataa_sig,
		AeB	 => AeB_sig,
		AgB	 => AgB_sig
	);

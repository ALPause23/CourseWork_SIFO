lpm_compare11_inst : lpm_compare11 PORT MAP (
		dataa	 => dataa_sig,
		AeB	 => AeB_sig
	);

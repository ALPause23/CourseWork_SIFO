lpm_bustri5_inst : lpm_bustri5 PORT MAP (
		data	 => data_sig,
		enabledt	 => enabledt_sig,
		tridata	 => tridata_sig
	);

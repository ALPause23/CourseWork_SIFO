lpm_compare1_inst : lpm_compare1 PORT MAP (
		dataa	 => dataa_sig,
		AgeB	 => AgeB_sig
	);

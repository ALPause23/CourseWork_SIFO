lpm_decode6_inst : lpm_decode6 PORT MAP (
		data	 => data_sig,
		enable	 => enable_sig,
		eq0	 => eq0_sig,
		eq1	 => eq1_sig,
		eq10	 => eq10_sig,
		eq11	 => eq11_sig,
		eq12	 => eq12_sig,
		eq13	 => eq13_sig,
		eq14	 => eq14_sig,
		eq15	 => eq15_sig,
		eq16	 => eq16_sig,
		eq17	 => eq17_sig,
		eq18	 => eq18_sig,
		eq19	 => eq19_sig,
		eq2	 => eq2_sig,
		eq20	 => eq20_sig,
		eq3	 => eq3_sig,
		eq4	 => eq4_sig,
		eq5	 => eq5_sig,
		eq6	 => eq6_sig,
		eq7	 => eq7_sig,
		eq8	 => eq8_sig,
		eq9	 => eq9_sig
	);

lpm_compare10_inst : lpm_compare10 PORT MAP (
		dataa	 => dataa_sig,
		AeB	 => AeB_sig,
		AlB	 => AlB_sig
	);

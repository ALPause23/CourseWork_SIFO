lpm_decode6_inst : lpm_decode6 PORT MAP (
		data	 => data_sig,
		eq1	 => eq1_sig,
		eq2	 => eq2_sig
	);

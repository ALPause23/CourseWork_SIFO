lpm_dff7_inst : lpm_dff7 PORT MAP (
		aload	 => aload_sig,
		clock	 => clock_sig,
		data	 => data_sig,
		q	 => q_sig
	);

lpm_compare5_inst : lpm_compare5 PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		AeB	 => AeB_sig
	);

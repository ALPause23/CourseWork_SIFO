lpm_counter5_inst : lpm_counter5 PORT MAP (
		aclr	 => aclr_sig,
		clock	 => clock_sig,
		sclr	 => sclr_sig,
		q	 => q_sig
	);

lpm_bustri2_inst : lpm_bustri2 PORT MAP (
		data	 => data_sig,
		enabledt	 => enabledt_sig,
		enabletr	 => enabletr_sig,
		result	 => result_sig,
		tridata	 => tridata_sig
	);

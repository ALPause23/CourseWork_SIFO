lpm_add_sub4_inst : lpm_add_sub4 PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		result	 => result_sig
	);

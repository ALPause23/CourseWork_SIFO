lpm_compare9_inst : lpm_compare9 PORT MAP (
		dataa	 => dataa_sig,
		AeB	 => AeB_sig
	);

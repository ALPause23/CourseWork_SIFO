lpm_compare6_inst : lpm_compare6 PORT MAP (
		dataa	 => dataa_sig,
		AeB	 => AeB_sig,
		AneB	 => AneB_sig
	);

lpm_compare12_inst : lpm_compare12 PORT MAP (
		dataa	 => dataa_sig,
		AeB	 => AeB_sig,
		AgB	 => AgB_sig,
		AlB	 => AlB_sig,
		AleB	 => AleB_sig
	);

lpm_compare13_inst : lpm_compare13 PORT MAP (
		dataa	 => dataa_sig,
		AeB	 => AeB_sig
	);

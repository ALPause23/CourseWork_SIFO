lpm_dff7_inst : lpm_dff7 PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		enable	 => enable_sig,
		q	 => q_sig
	);

lpm_compare7_inst : lpm_compare7 PORT MAP (
		dataa	 => dataa_sig,
		AeB	 => AeB_sig,
		AlB	 => AlB_sig
	);

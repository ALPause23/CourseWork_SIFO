lpm_counter2_inst : lpm_counter2 PORT MAP (
		clk_en	 => clk_en_sig,
		clock	 => clock_sig,
		sclr	 => sclr_sig,
		sset	 => sset_sig,
		cout	 => cout_sig,
		q	 => q_sig
	);

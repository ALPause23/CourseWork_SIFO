lpm_add_sub2_inst : lpm_add_sub2 PORT MAP (
		cin	 => cin_sig,
		dataa	 => dataa_sig,
		result	 => result_sig
	);

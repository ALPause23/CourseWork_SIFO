lpm_rom0_inst : lpm_rom0 PORT MAP (
		address	 => address_sig,
		inclock	 => inclock_sig,
		outclock	 => outclock_sig,
		q	 => q_sig
	);

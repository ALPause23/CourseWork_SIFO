lpm_compare8_inst : lpm_compare8 PORT MAP (
		dataa	 => dataa_sig,
		AeB	 => AeB_sig,
		AgB	 => AgB_sig,
		AleB	 => AleB_sig
	);

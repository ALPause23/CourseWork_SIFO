lpm_add_sub5_inst : lpm_add_sub5 PORT MAP (
		add_sub	 => add_sub_sig,
		dataa	 => dataa_sig,
		result	 => result_sig
	);
